package pkg;
    localparam WIDTH = 8;
    typedef logic [WIDTH-1:0]  data_t;
endpackage 