package afifo_tb_pkg;

localparam DW = 16;
typedef logic [DW-1] data_t;
typedef bit bit_t;

endpackage