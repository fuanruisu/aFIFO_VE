`ifndef MY_FIFO_PKTE
    `define FIFO_PKTE_SV
package afifo_pkg;

    localparam D_WIDTH = 8;
    typedef logic [D_WIDTH-1:0] data_ty;
    
endpackage
`endif