interface fifo(
    input clk
);